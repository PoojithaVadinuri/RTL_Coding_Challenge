
`include "top.sv"
`include "program.sv"


﻿
