module fa(s,cout,a,b,cin);

input a,b,cin;

output s,cout;

ha HA1(s1,c1,a,b);
ha HA2(s,c2,s1,cin);
or G1(cout,c1,c2);

endmodule