module fa(cout,sum,a,b,c);
input a,b,c;
output sum,cout;

ha h1(c0,s0,a,b);
ha h2(c1,sum,s0,c);
or h3(cout,c0,c1);
endmodule